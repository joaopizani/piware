process(sel, a, b)
begin
    if (sel = ‘0’) then
        y <= a;
    end if;
end process;
